module test_verilog()
//Register module instantition template. 
  //Will automate late.
endmodule 
